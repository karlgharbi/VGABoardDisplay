------------------------------------------------------------------------
-- mouse_displayer.vhd
------------------------------------------------------------------------
-- Author : Karl Gharbi
--          
------------------------------------------------------------------------
-- Software version : Xilinx ISE 7.1.04i
--                    WebPack
-- Device	        : 3s200ft256-4
------------------------------------------------------------------------
-- This file is a modification of the MouseDisplay sample code, designed by
-- Ulrich Zolt�n of Digilent. The goal is to have this file serve as a
-- generic flatbed to show game board graphics.
------------------------------------------------------------------------
--  Behavioral description
------------------------------------------------------------------------
-- Mouse position is received from the mouse_controller, horizontal and
-- vertical counters are received from vga_module and if the counters
-- are inside the mouse cursor bounds, then the mouse is sent to the
-- screen.
-- The mouse display module can be also used as an overlay of the VGA 
-- signal, also blanking the VGA screen, if the red_in, green_in, blue_in 
-- and the blank_in signals are used. 
-- In this application the signals mentioned and their corresponding code 
-- lines are commented, therefore the mouse display module only generates 
-- the RGB signals to display the cursor, and the VGA controller decides 
-- whether or not to display the cursor.
-- The mouse cursor is 16x16 pixels and uses 2 colors: white and black. 
-- For the color encoding 2 bits are used to be able to use transparency. 
-- The cursor is stored in a 256X2 bit distributed ram memory. If the current
-- pixel of the mouse is "00" then output color is black, if "01" then is
-- white and if "10" or "11" then the pixel is transparent and the input 
-- R, G and B signals are passed to the output. 
-- In this way, the mouse cursor will not be a 16x16 square, instead will 
-- have an arrow shape.
-- The memory address is composed from the difference of the vga counters
-- and mouse position: xdiff is the difference on 4 bits (because cursor
-- is 16 pixels width) between the horizontal vga counter and the xpos
-- of the mouse. ydiff is the difference on 4 bits (because cursor
-- has 16 pixels in height) between the vertical vga counter and the
-- ypos of the mouse. By concatenating ydiff and xidff (in this order)
-- the memory address of the current pixel is obtained.
-- A distributed memory implementation is forced by the attributes, to save 
-- BRAM resources.
-- If the blank input from the vga_module is active, this means that current
-- pixel is not inside visible screen and color outputs are set to black
------------------------------------------------------------------------
--  Port definitions
------------------------------------------------------------------------
-- pixel_clk      - input pin, representing the pixel clock, used
--                - by the vga_controller for the currently used
--                - resolution, generated by a dcm. 25MHz for 640x480,
--                - 40MHz for 800x600 and 108 MHz for 1280x1024. 
--                - This clock is used to read pixels from memory 
--                - and output data on color outputs.
-- hres           - input pin, 12 bits, from vga_module
--                - the horizontal resolution of the display to render to
--                - to be halved to center the board display.
-- vres           - input pin, 12 bits, from vga_module
--                - the vertical resolution of the display in question
--                - to be halved to center the board display.
-- hcount         - input pin, 12 bits, from vga_module
--                - the horizontal counter from the vga_controller
--                - tells the horizontal position of the current pixel
--                - on the screen from left to right.
-- vcount         - input pin, 12 bits, from vga_module
--                - the vertical counter from the vga_controller
--                - tells the vertical position of the currentl pixel
--                - on the screen from top to bottom.
-- red_out        - output pin, 4 bits, to vga hardware module.
--                - red output channel
-- green_out      - output pin, 4 bits, to vga hardware module.
--                - green output channel
-- blue_out       - output pin, 4 bits, to vga hardware module.
--                - blue output channel

------------------- Signals used when the mouse display is in overlay mode

-- blank          - input pin, from vga_module
--                - if active, current pixel is not in visible area,
--                - and color outputs should be set on 0.
-- red_in         - input pin, 4 bits, from effects_layer
--                - red channel input of the image to be displayed
-- green_in       - input pin, 4 bits, from effects_layer
--                - green channel input of the image to be displayed
-- blue_in        - input pin, 4 bits, from effects_layer
--                - blue channel input of the image to be displayed
------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.math_real.all;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.NUMERIC_STD.ALL;

-- simulation library
--library UNISIM;
--use UNISIM.VComponents.all;

-- the boardDisplay entity declaration
-- read above for behavioral description and port definitions.
entity BoardDisplay is
port (
   pixel_clk: in std_logic;

   hcount   : in std_logic_vector(11 downto 0);
   vcount   : in std_logic_vector(11 downto 0);
	
	hres     : in std_logic_vector(11 downto 0);
	vres     : in std_logic_vector(11 downto 0);
   --blank    : in std_logic; -- if VGA blank is used

   --red_in   : in std_logic_vector(3 downto 0); -- if VGA signal pass-through is used
   --green_in : in std_logic_vector(3 downto 0);
   --blue_in  : in std_logic_vector(3 downto 0);
   
   enable_display_out : out std_logic;

   red_out  : out std_logic_vector(3 downto 0);
   green_out: out std_logic_vector(3 downto 0);
   blue_out : out std_logic_vector(3 downto 0)
);

-- force synthesizer to extract distributed ram for the
-- displayrom signal, and not a block ram, to save BRAM resources.
attribute rom_extract : string;
attribute rom_extract of BoardDisplay: entity is "yes";
attribute rom_style : string;
attribute rom_style of BoardDisplay: entity is "distributed";

end BoardDisplay;

architecture Behavioral of BoardDisplay is

------------------------------------------------------------------------
-- CONSTANTS
------------------------------------------------------------------------

constant numRows: integer := 6;
constant numColumns: integer := 7;
constant slotSize: integer := 100;
constant borderSize: integer := 10;

constant displayWidth: integer := ((numColumns * slotSize) + ((numColumns+1) * borderSize));
constant displayHeight: integer := (((numRows+1 * slotSize) + ((numRows+1) * borderSize) + borderSize));

constant X_OFFSET: std_logic_vector(11 downto 0) := std_logic_vector(to_unsigned(displayHeight, 12));
constant Y_OFFSET: std_logic_vector(11 downto 0) := std_logic_vector(to_unsigned(displayWidth, 12));
						
constant X_OFFSET_HALF: std_logic_vector(11 downto 0) := '0' & X_OFFSET(11 downto 1);
constant Y_OFFSET_HALF: std_logic_vector(11 downto 0) := '0' & Y_OFFSET(11 downto 1);

type newColumn is array (displayWidth downto 0) of std_logic_vector(1 downto 0);
--change: Use 3D array rather than 2D array in order to accommodate rectangular spritemap
type newdisplayram is array (displayHeight downto 0) of newColumn;
type displayRom is array(0 to 28, 43 downto 0) of std_logic_vector(1 downto 0);
-- the memory that holds the cursor.
-- change: 00 now represents transparent instead of black (i dun goofed)
-- change: I take that back
-- 00 - black
-- 01 - yellow
-- 1x - transparent

constant board: displayrom := (

("01","01","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","01","01"),
("01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01"),
("01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01"),
("01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01"),
("01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01"),
("01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01"),
("01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01"),
("01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01"),
("01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01"),
("01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01"),
("01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01"),
("01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01"),
("01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01"),
("01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01"),
("01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01"),
("01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01"),
("01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01"),
("01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01"),
("01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01"),
("01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01"),
("01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01"),
("01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01"),
("01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01"),
("01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01"),
("01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01","00","00","00","00","00","01","01"),
("01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01"),
("01","01","01","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","01","01","01"),
("01","01","01","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","01","01","01"),
("01","01","01","01","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","01","01","01","01")

);

-- width and height of cursor.
-- change: Use seperate offsets for horizontal and vertical dimensions
--constant X_OFFSET: std_logic_vector(5 downto 0) := "101100";   -- 44
--constant Y_OFFSET: std_logic_vector(4 downto 0) := "11101"; --29
--
--constant X_OFFSET_HALF: std_logic_vector(4 downto 0) := X_OFFSET(5 downto 1);
--constant Y_OFFSET_HALF: std_logic_vector(3 downto 0) := Y_OFFSET(4 downto 1);

--44x28 bitmap, not square
--Will determine how to properly express this
--When picking the differential, will need to limit the max value to be
--within the space of the actual ROM
--(2^6 + 2^5 = 11 bits for ROM address)
--2048 values max for 11 bit number
--1276 addresses used

------------------------------------------------------------------------
-- SIGNALS
------------------------------------------------------------------------
--new: provide information for where the top left corner of the board will be,
--as mouse input will not be used to figure that out.
--coded as signals, but in practice considered to be a constant.
signal hPoint : std_logic_vector(11 downto 0) := ('0' & hres(11 downto 1)) + X_OFFSET_HALF;
signal vPoint : std_logic_vector(11 downto 0) := ('0' & vres(11 downto 1)) + Y_OFFSET_HALF;

--newer: New board replacement code
signal newBoard : newdisplayram;
signal boardMade : std_logic := '0';

-- pixel from the display memory, representing currently displayed
-- pixel of the cursor, if the cursor is being display at this point
signal boardpixel: std_logic_vector(1 downto 0) := (others => '0');
-- when high, enables displaying of the cursor, and reading the
-- cursor memory.
signal enable_display: std_logic := '0';

-- difference in range 0-15 between the vga counters and mouse position
--change: xdiff and ydiff lengths, per bitmap change
--signal xdiff: std_logic_vector(5 downto 0) := (others => '0');
--signal ydiff: std_logic_vector(4 downto 0) := (others => '0');
signal xdiff: std_logic_vector(11 downto 0) := (others => '0');
signal ydiff: std_logic_vector(11 downto 0) := (others => '0');

signal red_int  : std_logic_vector(3 downto 0);
signal green_int: std_logic_vector(3 downto 0);
signal blue_int : std_logic_vector(3 downto 0);

signal red_int1  : std_logic_vector(3 downto 0);
signal green_int1: std_logic_vector(3 downto 0);
signal blue_int1 : std_logic_vector(3 downto 0);

begin

--what did I want to do
--Board size has been determined, based on predetermined # of lines & thickness
--For each row, have (x+1) divisions and x slots, where x is the number of slots
--Except for the first row, which will only have divisions at the ends.
--So, what shall the structure be?
--Initial loop: For (slot height), fill (borderSize) at beginning and end, rest is blank
--Main loop: For(slot height * rowCount), fill with (borderSize), then blank for slotSize, repeat 
--until (x+1) divisions done
--Final Loop: Generate legs
--	--generate/update new board
	makeBoard: process(pixel_clk, newBoard, boardMade)
	begin
		if(boardMade = '0') then
			for row in 0 to displayWidth loop
				for column in 0 to displayHeight loop
					--top part generation conditionals
					if(row < (slotSize)) then
						if((column < borderSize) or (column > (X_OFFSET - 1 - borderSize))) then
							newBoard(row(column)) <= "01";
						else
							newBoard(row(column)) <= "00";
						end if;
				   --bottom part generation conditionals
					elsif(row >= ((numRows+1) * (borderSize + slotSize))) then
						if((column < (Y_OFFSET - (numRows+1) * (borderSize + slotSize))) or
							(column > (Y_OFFSET - (Y_OFFSET - (numRows+1) * (borderSize + slotSize))))) then
							newBoard(row, column) <= "01";
						else
							newBoard(row, column) <= "00";
						end if;
					--main board generation conditionals
					else
						--slot row generation conditionals
						if((row mod (slotSize + borderSize)) < slotSize) then
							if((column mod (slotSize + borderSize)) < borderSize) then
								newBoard(row, column) <= "01";
							else
								newBoard(row, column) <= "00";
							end if;
						--border row generation conditional
						else
							newBoard(row) <= (others => "01");
						end if;
					end if;
				end loop;
			end loop;
		boardMade <= '1';
		end if;
	end process;
		

--   -- compute xdiff
--   x_diff: process(hcount, hPoint)
--   variable temp_diff: std_logic_vector(11 downto 0) := (others => '0');
--   begin
--			temp_diff := hcount - hPoint;
--			if (temp_diff(5 downto 0) > X"2B") then --X"2B" = 43
--				xdiff <= "101011";
--			else
--				xdiff <= temp_diff(5 downto 0);
--			end if;
--   end process x_diff;
--
--   -- compute ydiff
--   y_diff: process(vcount, vPoint)
--   variable temp_diff: std_logic_vector(11 downto 0) := (others => '0');
--   begin
--         temp_diff := vcount - vPoint;
--			if (temp_diff(4 downto 0) > X"1C") then --X"1C" = 28
--				ydiff <= "11100";
--			else
--				ydiff <= temp_diff(4 downto 0);
--			end if;
--   end process y_diff;

-- compute xdiff
	x_diff: process(hcount, hPoint)
   variable temp_diff: std_logic_vector(11 downto 0) := (others => '0');
   begin
			temp_diff := hcount - hPoint;
			if (temp_diff > X_OFFSET) then
				xdiff <= X_OFFSET;
			else
				xdiff <= temp_diff;
			end if;
   end process x_diff;
	
	   -- compute ydiff
   y_diff: process(vcount, vPoint)
   variable temp_diff: std_logic_vector(11 downto 0) := (others => '0');
   begin
         temp_diff := vcount - vPoint;
			if (temp_diff > Y_OFFSET) then --X"1C" = 28
				ydiff <= Y_OFFSET;
			else
				ydiff <= temp_diff;
			end if;
   end process y_diff;

 -- read pixel from memory at address obtained by concatenation of
   -- ydiff and xdiff
--	boardpixel <= board(conv_integer(ydiff), conv_integer(xdiff))
--                 when rising_edge(pixel_clk);
   boardpixel <= newBoard(conv_integer(ydiff), conv_integer(xdiff))
                 when rising_edge(pixel_clk);

   -- set enable_mouse_display high if vga counters inside cursor block
	--change: OFFSET replaced with X_OFFSET and Y_OFFSET for hcount and vcount
   enable_display_control: process(pixel_clk, hcount, vcount, hPoint, vPoint)
   begin
      if(rising_edge(pixel_clk)) then
         if(hcount >= hPoint + 1 and hcount <= (hPoint + X_OFFSET) and
            vcount >= vPoint + 1 and vcount <= (vPoint + Y_OFFSET)) and
            (boardpixel = "01" or boardpixel = "00")
         then
            enable_display <= '1';
         else
            enable_display <= '0';
         end if;
      end if;
   end process enable_display_control;
   
enable_display_out <= enable_display;

   -- if cursor display is enabled, then, according to pixel
   -- value, set the output color channels.
 process(pixel_clk)
   begin
      if(rising_edge(pixel_clk)) then
         -- if in visible screen
--       if(blank = '0') then
            -- in display is enabled
            if(enable_display = '1') then
               -- yellow pixel of cursor
					--change: white -> yellow
               if(boardpixel = "01") then
                  red_out <= (others => '1');
                  green_out <= (others => '1');
                  blue_out <= (others => '0');
               -- black pixel of cursor
               elsif(boardpixel = "00") then
                  red_out <= (others => '0');
                  green_out <= (others => '0');
                  blue_out <= (others => '0');
               -- transparent pixel of cursor
               -- let input pass to output
--               else
--                  red_out <= red_in;
--                  green_out <= green_in;
--                  blue_out <= blue_in;
               end if;
            -- cursor display is not enabled
            -- let input pass to output.
--          else
--               red_out <= red_in;
--               green_out <= green_in;
--               blue_out <= blue_in;
            end if;
         -- not in visible screen, black outputs.
--       else
--            red_out <= (others => '0');
--            green_out <= (others => '0');
--            blue_out <= (others => '0');
--      end if;
      end if;
   end process;


end Behavioral;
